`timescale 1ns / 1ps
//------------------------------------------------------------------------------
// Release Date  : 25_07_2022
// Design Name   : FPGA CLB Resources
// Release       : 0.3 
// Module Name   : mux_16to1.v
// Target Devices: Xilinx 7 series FPGA
// Tool versions : VIVADO 2020.1
// Description   : 16 to 1 Multiplexer		   
//------------------------------------------------------------------------------
// DESIGN HIERARCHY 
// - No - Basic Module
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
// MODULE DECLARATION 
//------------------------------------------------------------------------------  
  module mux_16to1 
  (
//------------------------------------------------------------------------------
// INPUT DECLARATION
//------------------------------------------------------------------------------ 
    input [ 15:0] mux_inp	,	// multiplex inputs declaration   
    input [  3:0]     sel	,	// select inputs declaration
//------------------------------------------------------------------------------
// OUTPUT DECLARATION
//------------------------------------------------------------------------------
    output 	 mux_out		// multiplex output declaration 
  ); 
//------------------------------------------------------------------------------
// DATAFLOW MODELING - MUX LOGIC
//------------------------------------------------------------------------------
  assign mux_out = mux_inp[sel] ;   

endmodule 
