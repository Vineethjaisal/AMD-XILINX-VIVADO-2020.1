`timescale 1ns / 1ps
//------------------------------------------------------------------------------
// Release Date  : 25_07_2022
// Design Name   : FPGA CLB Resources
// Release       : 0.3 
// Module Name   : adder_8bit.v
// Target Devices: Xilinx 7 series FPGA
// Tool versions : VIVADO 2020.1
// Description   : 8 bit Adder		   
//------------------------------------------------------------------------------
// DESIGN HIERARCHY 
// - No - Basic Module
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
// MODULE DECLARATION 
//------------------------------------------------------------------------------  
  module adder_8bit 
  (
//------------------------------------------------------------------------------
// INPUT DECLARATION
//------------------------------------------------------------------------------ 
    input 	[7:0]		a	,	// input a declaration 
    input 	[7:0]		b	,	// input b declaration
//------------------------------------------------------------------------------
// OUTPUT DECLARATION
//------------------------------------------------------------------------------
    output 	[8:0]		sum		// output full adder sum declaration 
  ); 
//------------------------------------------------------------------------------
// DATA FLOW MODELING - ADDTION LOGIC
//------------------------------------------------------------------------------
  assign sum  =  a + b 	;
  
endmodule 
