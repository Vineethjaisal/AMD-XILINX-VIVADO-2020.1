`timescale 1ns / 1ps
//------------------------------------------------------------------------------
// Release Date  : 25_07_2022
// Design Name   : FPGA CLB Resources
// Release       : 0.3 
// Module Name   : sp_dist_ram_256x8.v
// Target Devices: Xilinx 7 series FPGA
// Tool versions : VIVADO 2020.1
// Description   : Single Port RAM Asynchronous Read - Distributed RAM		   
//------------------------------------------------------------------------------
// DESIGN HIERARCHY 
// - No - Basic Module
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
// MODULE DECLARATION 
//------------------------------------------------------------------------------
  module sp_dist_ram_256x8
  (
//------------------------------------------------------------------------------
// INPUT DECLARATION
//------------------------------------------------------------------------------
  input 	    clk_in		     		, // Clock Input
  input         write_en			, // Write Enable Logic
  input  [7:0]  address_in	     		, // 8 bit Address Bus
  input  [7:0]  data_in				, // 8 bit Input Data Bus 
//------------------------------------------------------------------------------
// OUTPUT DECLARATION
//------------------------------------------------------------------------------
  output [7:0]	data_out	  	          // 8 bit Output Data Bus
  ); 
//------------------------------------------------------------------------------
// MEMORY ARRAY DECLARATION
//------------------------------------------------------------------------------
  reg 	 [7:0]  dram_mem [0:255]  		; // RAM Memory Array 
//------------------------------------------------------------------------------
//[7][6][5][4][3][2][1][0] - 0
//[7][6][5][4][3][2][1][0] - 1
//[7][6][5][4][3][2][1][0] - 2
//[0][0][0][0][0][1][0][1] - 3 //data_in = 5
//[7][6][5][4][3][2][1][0] - 4
//[7][6][5][4][3][2][1][0] - 5
//[7][6][5][4][3][2][1][0] - 6
//------------------------
//------------------------
//------------------------
//[7][6][5][4][3][2][1][0] - 252
//[7][6][5][4][3][2][1][0] - 253
//[7][6][5][4][3][2][1][0] - 254
//[7][6][5][4][3][2][1][0] - 255
//------------------------------------------------------------------------------
// PROCEDURAL ALWAYS BLOCK - Distributed RAM Write / Read Logic 
//------------------------------------------------------------------------------     
  always@(posedge clk_in)
    begin
      if(write_en)
         begin
           dram_mem[address_in] <= data_in	; // Sync. Write  
         end
    end


  assign data_out = dram_mem[address_in]  	; // Async. Read  

endmodule
